`include "c17.v"
module c17_tb;
reg N1;
reg N2;
reg N3;
reg N6;
reg N7;

wire N22;
wire N23;

initial begin
	$dumpfile("c17_tb.vcd");
	$dumpvars(0, c17_tb);
	$monitor($time, ": , N1: %b(%d), N2: %b(%d), N3: %b(%d), N6: %b(%d), N7: %b(%d), N22: %b(%d), N23: %b(%d)", N1, N1, N2, N2, N3, N3, N6, N6, N7, N7, N22, N22, N23, N23);
end
c17 c17_(.N1(N1), .N2(N2), .N3(N3), .N6(N6), .N7(N7), .N22(N22), .N23(N23));


initial begin
N1 = 1'b0; 
N2 = 1'b0; 
N3 = 1'b0; 
N6 = 1'b0; 
N7 = 1'b0; 

#10 N1 = 1'b1; N2 = 1'b0; N3 = 1'b0; N6 = 1'b0; N7 = 1'b0; 
#10 N1 = 1'b0; N2 = 1'b1; N3 = 1'b0; N6 = 1'b0; N7 = 1'b0; 
#10 N1 = 1'b1; N2 = 1'b1; N3 = 1'b0; N6 = 1'b0; N7 = 1'b0; 
#10 N1 = 1'b0; N2 = 1'b0; N3 = 1'b1; N6 = 1'b0; N7 = 1'b0; 
#10 N1 = 1'b1; N2 = 1'b0; N3 = 1'b1; N6 = 1'b0; N7 = 1'b0; 
#10 N1 = 1'b0; N2 = 1'b1; N3 = 1'b1; N6 = 1'b0; N7 = 1'b0; 
#10 N1 = 1'b1; N2 = 1'b1; N3 = 1'b1; N6 = 1'b0; N7 = 1'b0; 
#10 N1 = 1'b0; N2 = 1'b0; N3 = 1'b0; N6 = 1'b1; N7 = 1'b0; 
#10 N1 = 1'b1; N2 = 1'b0; N3 = 1'b0; N6 = 1'b1; N7 = 1'b0; 
#10 N1 = 1'b0; N2 = 1'b1; N3 = 1'b0; N6 = 1'b1; N7 = 1'b0; 
#10 N1 = 1'b1; N2 = 1'b1; N3 = 1'b0; N6 = 1'b1; N7 = 1'b0; 
#10 N1 = 1'b0; N2 = 1'b0; N3 = 1'b1; N6 = 1'b1; N7 = 1'b0; 
#10 N1 = 1'b1; N2 = 1'b0; N3 = 1'b1; N6 = 1'b1; N7 = 1'b0; 
#10 N1 = 1'b0; N2 = 1'b1; N3 = 1'b1; N6 = 1'b1; N7 = 1'b0; 
#10 N1 = 1'b1; N2 = 1'b1; N3 = 1'b1; N6 = 1'b1; N7 = 1'b0; 
#10 N1 = 1'b0; N2 = 1'b0; N3 = 1'b0; N6 = 1'b0; N7 = 1'b1; 
#10 N1 = 1'b1; N2 = 1'b0; N3 = 1'b0; N6 = 1'b0; N7 = 1'b1; 
#10 N1 = 1'b0; N2 = 1'b1; N3 = 1'b0; N6 = 1'b0; N7 = 1'b1; 
#10 N1 = 1'b1; N2 = 1'b1; N3 = 1'b0; N6 = 1'b0; N7 = 1'b1; 
#10 N1 = 1'b0; N2 = 1'b0; N3 = 1'b1; N6 = 1'b0; N7 = 1'b1; 
#10 N1 = 1'b1; N2 = 1'b0; N3 = 1'b1; N6 = 1'b0; N7 = 1'b1; 
#10 N1 = 1'b0; N2 = 1'b1; N3 = 1'b1; N6 = 1'b0; N7 = 1'b1; 
#10 N1 = 1'b1; N2 = 1'b1; N3 = 1'b1; N6 = 1'b0; N7 = 1'b1; 
#10 N1 = 1'b0; N2 = 1'b0; N3 = 1'b0; N6 = 1'b1; N7 = 1'b1; 
#10 N1 = 1'b1; N2 = 1'b0; N3 = 1'b0; N6 = 1'b1; N7 = 1'b1; 
#10 N1 = 1'b0; N2 = 1'b1; N3 = 1'b0; N6 = 1'b1; N7 = 1'b1; 
#10 N1 = 1'b1; N2 = 1'b1; N3 = 1'b0; N6 = 1'b1; N7 = 1'b1; 
#10 N1 = 1'b0; N2 = 1'b0; N3 = 1'b1; N6 = 1'b1; N7 = 1'b1; 
#10 N1 = 1'b1; N2 = 1'b0; N3 = 1'b1; N6 = 1'b1; N7 = 1'b1; 
#10 N1 = 1'b0; N2 = 1'b1; N3 = 1'b1; N6 = 1'b1; N7 = 1'b1; 
#10 N1 = 1'b1; N2 = 1'b1; N3 = 1'b1; N6 = 1'b1; N7 = 1'b1; 
#10 N1 = 1'b0; N2 = 1'b0; N3 = 1'b0; N6 = 1'b0; N7 = 1'b0; 

end
endmodule
