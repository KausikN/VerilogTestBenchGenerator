`include "c432.v"
module c432_tb;
reg N1;
reg N4;
reg N8;
reg N11;
reg N14;
reg N17;
reg N21;
reg N24;
reg N27;
reg N30;
reg N34;
reg N37;
reg N40;
reg N43;
reg N47;
reg N50;
reg N53;
reg N56;
reg N60;
reg N63;
reg N66;
reg N69;
reg N73;
reg N76;
reg N79;
reg N82;
reg N86;
reg N89;
reg N92;
reg N95;
reg N99;
reg N102;
reg N105;
reg N108;
reg N112;
reg N115;

wire N223;
wire N329;
wire N370;
wire N421;
wire N430;
wire N431;
wire N432;

initial begin
	$dumpfile("c432_tb.vcd");
	$dumpvars(0, c432_tb);
	$monitor($time, ": , N1: %b(%d), N4: %b(%d), N8: %b(%d), N11: %b(%d), N14: %b(%d), N17: %b(%d), N21: %b(%d), N24: %b(%d), N27: %b(%d), N30: %b(%d), N34: %b(%d), N37: %b(%d), N40: %b(%d), N43: %b(%d), N47: %b(%d), N50: %b(%d), N53: %b(%d), N56: %b(%d), N60: %b(%d), N63: %b(%d), N66: %b(%d), N69: %b(%d), N73: %b(%d), N76: %b(%d), N79: %b(%d), N82: %b(%d), N86: %b(%d), N89: %b(%d), N92: %b(%d), N95: %b(%d), N99: %b(%d), N102: %b(%d), N105: %b(%d), N108: %b(%d), N112: %b(%d), N115: %b(%d), N223: %b(%d), N329: %b(%d), N370: %b(%d), N421: %b(%d), N430: %b(%d), N431: %b(%d), N432: %b(%d)", N1, N1, N4, N4, N8, N8, N11, N11, N14, N14, N17, N17, N21, N21, N24, N24, N27, N27, N30, N30, N34, N34, N37, N37, N40, N40, N43, N43, N47, N47, N50, N50, N53, N53, N56, N56, N60, N60, N63, N63, N66, N66, N69, N69, N73, N73, N76, N76, N79, N79, N82, N82, N86, N86, N89, N89, N92, N92, N95, N95, N99, N99, N102, N102, N105, N105, N108, N108, N112, N112, N115, N115, N223, N223, N329, N329, N370, N370, N421, N421, N430, N430, N431, N431, N432, N432);
end
c432 c432_(.N1(N1), .N4(N4), .N8(N8), .N11(N11), .N14(N14), .N17(N17), .N21(N21), .N24(N24), .N27(N27), .N30(N30), .N34(N34), .N37(N37), .N40(N40), .N43(N43), .N47(N47), .N50(N50), .N53(N53), .N56(N56), .N60(N60), .N63(N63), .N66(N66), .N69(N69), .N73(N73), .N76(N76), .N79(N79), .N82(N82), .N86(N86), .N89(N89), .N92(N92), .N95(N95), .N99(N99), .N102(N102), .N105(N105), .N108(N108), .N112(N112), .N115(N115), .N223(N223), .N329(N329), .N370(N370), .N421(N421), .N430(N430), .N431(N431), .N432(N432));


initial begin
N1 = 1'b0; 
N4 = 1'b0; 
N8 = 1'b0; 
N11 = 1'b0; 
N14 = 1'b0; 
N17 = 1'b0; 
N21 = 1'b0; 
N24 = 1'b0; 
N27 = 1'b0; 
N30 = 1'b0; 
N34 = 1'b0; 
N37 = 1'b0; 
N40 = 1'b0; 
N43 = 1'b0; 
N47 = 1'b0; 
N50 = 1'b0; 
N53 = 1'b0; 
N56 = 1'b0; 
N60 = 1'b0; 
N63 = 1'b0; 
N66 = 1'b0; 
N69 = 1'b0; 
N73 = 1'b0; 
N76 = 1'b0; 
N79 = 1'b0; 
N82 = 1'b0; 
N86 = 1'b0; 
N89 = 1'b0; 
N92 = 1'b0; 
N95 = 1'b0; 
N99 = 1'b0; 
N102 = 1'b0; 
N105 = 1'b0; 
N108 = 1'b0; 
N112 = 1'b0; 
N115 = 1'b0; 

#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b0; N11 = 1'b0; N14 = 1'b0; N17 = 1'b1; N21 = 1'b1; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b0; N37 = 1'b0; N40 = 1'b0; N43 = 1'b0; N47 = 1'b1; N50 = 1'b0; N53 = 1'b1; N56 = 1'b1; N60 = 1'b1; N63 = 1'b0; N66 = 1'b1; N69 = 1'b1; N73 = 1'b1; N76 = 1'b0; N79 = 1'b0; N82 = 1'b1; N86 = 1'b1; N89 = 1'b0; N92 = 1'b0; N95 = 1'b0; N99 = 1'b1; N102 = 1'b0; N105 = 1'b1; N108 = 1'b1; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b1; N11 = 1'b0; N14 = 1'b1; N17 = 1'b1; N21 = 1'b1; N24 = 1'b1; N27 = 1'b0; N30 = 1'b0; N34 = 1'b0; N37 = 1'b0; N40 = 1'b1; N43 = 1'b0; N47 = 1'b0; N50 = 1'b0; N53 = 1'b0; N56 = 1'b1; N60 = 1'b1; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b0; N76 = 1'b1; N79 = 1'b1; N82 = 1'b0; N86 = 1'b0; N89 = 1'b0; N92 = 1'b1; N95 = 1'b0; N99 = 1'b1; N102 = 1'b0; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b0; N11 = 1'b0; N14 = 1'b1; N17 = 1'b0; N21 = 1'b0; N24 = 1'b1; N27 = 1'b1; N30 = 1'b0; N34 = 1'b1; N37 = 1'b0; N40 = 1'b1; N43 = 1'b0; N47 = 1'b1; N50 = 1'b0; N53 = 1'b0; N56 = 1'b0; N60 = 1'b0; N63 = 1'b0; N66 = 1'b1; N69 = 1'b0; N73 = 1'b0; N76 = 1'b0; N79 = 1'b0; N82 = 1'b1; N86 = 1'b0; N89 = 1'b1; N92 = 1'b0; N95 = 1'b1; N99 = 1'b1; N102 = 1'b0; N105 = 1'b1; N108 = 1'b1; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b0; N11 = 1'b0; N14 = 1'b0; N17 = 1'b0; N21 = 1'b0; N24 = 1'b0; N27 = 1'b0; N30 = 1'b1; N34 = 1'b0; N37 = 1'b1; N40 = 1'b1; N43 = 1'b0; N47 = 1'b0; N50 = 1'b1; N53 = 1'b0; N56 = 1'b0; N60 = 1'b0; N63 = 1'b0; N66 = 1'b1; N69 = 1'b0; N73 = 1'b1; N76 = 1'b1; N79 = 1'b1; N82 = 1'b1; N86 = 1'b1; N89 = 1'b1; N92 = 1'b1; N95 = 1'b0; N99 = 1'b1; N102 = 1'b1; N105 = 1'b0; N108 = 1'b1; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b0; N11 = 1'b1; N14 = 1'b1; N17 = 1'b1; N21 = 1'b1; N24 = 1'b0; N27 = 1'b0; N30 = 1'b0; N34 = 1'b1; N37 = 1'b0; N40 = 1'b1; N43 = 1'b1; N47 = 1'b0; N50 = 1'b0; N53 = 1'b0; N56 = 1'b1; N60 = 1'b0; N63 = 1'b1; N66 = 1'b0; N69 = 1'b0; N73 = 1'b0; N76 = 1'b1; N79 = 1'b0; N82 = 1'b1; N86 = 1'b1; N89 = 1'b0; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b1; N105 = 1'b1; N108 = 1'b0; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b1; N11 = 1'b1; N14 = 1'b1; N17 = 1'b1; N21 = 1'b0; N24 = 1'b0; N27 = 1'b0; N30 = 1'b0; N34 = 1'b0; N37 = 1'b1; N40 = 1'b0; N43 = 1'b0; N47 = 1'b1; N50 = 1'b0; N53 = 1'b1; N56 = 1'b1; N60 = 1'b1; N63 = 1'b0; N66 = 1'b1; N69 = 1'b0; N73 = 1'b1; N76 = 1'b0; N79 = 1'b0; N82 = 1'b1; N86 = 1'b1; N89 = 1'b0; N92 = 1'b1; N95 = 1'b1; N99 = 1'b0; N102 = 1'b1; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b0; N8 = 1'b0; N11 = 1'b0; N14 = 1'b0; N17 = 1'b0; N21 = 1'b0; N24 = 1'b0; N27 = 1'b0; N30 = 1'b0; N34 = 1'b0; N37 = 1'b1; N40 = 1'b0; N43 = 1'b1; N47 = 1'b0; N50 = 1'b1; N53 = 1'b0; N56 = 1'b0; N60 = 1'b1; N63 = 1'b0; N66 = 1'b0; N69 = 1'b0; N73 = 1'b0; N76 = 1'b0; N79 = 1'b1; N82 = 1'b0; N86 = 1'b1; N89 = 1'b1; N92 = 1'b0; N95 = 1'b0; N99 = 1'b1; N102 = 1'b0; N105 = 1'b1; N108 = 1'b1; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b1; N11 = 1'b1; N14 = 1'b0; N17 = 1'b0; N21 = 1'b1; N24 = 1'b1; N27 = 1'b0; N30 = 1'b1; N34 = 1'b0; N37 = 1'b1; N40 = 1'b1; N43 = 1'b0; N47 = 1'b0; N50 = 1'b0; N53 = 1'b1; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b0; N69 = 1'b0; N73 = 1'b1; N76 = 1'b0; N79 = 1'b1; N82 = 1'b0; N86 = 1'b0; N89 = 1'b0; N92 = 1'b1; N95 = 1'b0; N99 = 1'b1; N102 = 1'b0; N105 = 1'b1; N108 = 1'b0; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b0; N8 = 1'b0; N11 = 1'b1; N14 = 1'b1; N17 = 1'b0; N21 = 1'b1; N24 = 1'b1; N27 = 1'b0; N30 = 1'b0; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b1; N47 = 1'b0; N50 = 1'b0; N53 = 1'b1; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b1; N69 = 1'b1; N73 = 1'b1; N76 = 1'b0; N79 = 1'b0; N82 = 1'b0; N86 = 1'b0; N89 = 1'b0; N92 = 1'b1; N95 = 1'b1; N99 = 1'b1; N102 = 1'b1; N105 = 1'b1; N108 = 1'b0; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b0; N11 = 1'b1; N14 = 1'b1; N17 = 1'b0; N21 = 1'b0; N24 = 1'b1; N27 = 1'b1; N30 = 1'b0; N34 = 1'b0; N37 = 1'b1; N40 = 1'b1; N43 = 1'b0; N47 = 1'b1; N50 = 1'b0; N53 = 1'b1; N56 = 1'b1; N60 = 1'b0; N63 = 1'b1; N66 = 1'b1; N69 = 1'b0; N73 = 1'b0; N76 = 1'b1; N79 = 1'b1; N82 = 1'b0; N86 = 1'b0; N89 = 1'b0; N92 = 1'b1; N95 = 1'b0; N99 = 1'b0; N102 = 1'b0; N105 = 1'b0; N108 = 1'b1; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b0; N11 = 1'b0; N14 = 1'b1; N17 = 1'b0; N21 = 1'b1; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b0; N37 = 1'b0; N40 = 1'b1; N43 = 1'b1; N47 = 1'b1; N50 = 1'b1; N53 = 1'b0; N56 = 1'b0; N60 = 1'b0; N63 = 1'b0; N66 = 1'b0; N69 = 1'b0; N73 = 1'b1; N76 = 1'b1; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b0; N92 = 1'b0; N95 = 1'b0; N99 = 1'b1; N102 = 1'b0; N105 = 1'b1; N108 = 1'b1; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b0; N11 = 1'b1; N14 = 1'b1; N17 = 1'b1; N21 = 1'b1; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b1; N37 = 1'b0; N40 = 1'b1; N43 = 1'b1; N47 = 1'b0; N50 = 1'b1; N53 = 1'b1; N56 = 1'b1; N60 = 1'b1; N63 = 1'b1; N66 = 1'b1; N69 = 1'b1; N73 = 1'b0; N76 = 1'b1; N79 = 1'b0; N82 = 1'b1; N86 = 1'b1; N89 = 1'b0; N92 = 1'b0; N95 = 1'b0; N99 = 1'b1; N102 = 1'b1; N105 = 1'b1; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b0; N8 = 1'b1; N11 = 1'b0; N14 = 1'b0; N17 = 1'b0; N21 = 1'b1; N24 = 1'b1; N27 = 1'b1; N30 = 1'b0; N34 = 1'b1; N37 = 1'b1; N40 = 1'b1; N43 = 1'b0; N47 = 1'b1; N50 = 1'b0; N53 = 1'b0; N56 = 1'b0; N60 = 1'b0; N63 = 1'b1; N66 = 1'b0; N69 = 1'b1; N73 = 1'b0; N76 = 1'b0; N79 = 1'b1; N82 = 1'b1; N86 = 1'b1; N89 = 1'b1; N92 = 1'b1; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b0; N108 = 1'b1; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b1; N11 = 1'b1; N14 = 1'b0; N17 = 1'b1; N21 = 1'b1; N24 = 1'b1; N27 = 1'b1; N30 = 1'b1; N34 = 1'b0; N37 = 1'b1; N40 = 1'b0; N43 = 1'b1; N47 = 1'b1; N50 = 1'b0; N53 = 1'b0; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b1; N76 = 1'b1; N79 = 1'b1; N82 = 1'b1; N86 = 1'b1; N89 = 1'b1; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b1; N108 = 1'b0; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b0; N8 = 1'b1; N11 = 1'b0; N14 = 1'b0; N17 = 1'b0; N21 = 1'b1; N24 = 1'b0; N27 = 1'b0; N30 = 1'b0; N34 = 1'b0; N37 = 1'b0; N40 = 1'b0; N43 = 1'b0; N47 = 1'b0; N50 = 1'b0; N53 = 1'b1; N56 = 1'b0; N60 = 1'b1; N63 = 1'b0; N66 = 1'b0; N69 = 1'b0; N73 = 1'b0; N76 = 1'b1; N79 = 1'b1; N82 = 1'b1; N86 = 1'b1; N89 = 1'b1; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b1; N105 = 1'b0; N108 = 1'b1; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b0; N8 = 1'b1; N11 = 1'b0; N14 = 1'b1; N17 = 1'b1; N21 = 1'b0; N24 = 1'b1; N27 = 1'b1; N30 = 1'b1; N34 = 1'b0; N37 = 1'b1; N40 = 1'b0; N43 = 1'b0; N47 = 1'b1; N50 = 1'b1; N53 = 1'b0; N56 = 1'b0; N60 = 1'b1; N63 = 1'b1; N66 = 1'b1; N69 = 1'b1; N73 = 1'b1; N76 = 1'b1; N79 = 1'b0; N82 = 1'b1; N86 = 1'b1; N89 = 1'b0; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b1; N108 = 1'b1; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b1; N11 = 1'b1; N14 = 1'b1; N17 = 1'b1; N21 = 1'b0; N24 = 1'b1; N27 = 1'b0; N30 = 1'b1; N34 = 1'b1; N37 = 1'b1; N40 = 1'b1; N43 = 1'b1; N47 = 1'b0; N50 = 1'b1; N53 = 1'b1; N56 = 1'b1; N60 = 1'b1; N63 = 1'b1; N66 = 1'b1; N69 = 1'b1; N73 = 1'b0; N76 = 1'b0; N79 = 1'b0; N82 = 1'b1; N86 = 1'b1; N89 = 1'b1; N92 = 1'b1; N95 = 1'b0; N99 = 1'b1; N102 = 1'b0; N105 = 1'b1; N108 = 1'b1; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b1; N11 = 1'b0; N14 = 1'b1; N17 = 1'b0; N21 = 1'b1; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b1; N37 = 1'b0; N40 = 1'b1; N43 = 1'b1; N47 = 1'b0; N50 = 1'b1; N53 = 1'b0; N56 = 1'b0; N60 = 1'b1; N63 = 1'b0; N66 = 1'b1; N69 = 1'b1; N73 = 1'b1; N76 = 1'b0; N79 = 1'b1; N82 = 1'b0; N86 = 1'b1; N89 = 1'b0; N92 = 1'b0; N95 = 1'b0; N99 = 1'b1; N102 = 1'b1; N105 = 1'b0; N108 = 1'b1; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b1; N11 = 1'b0; N14 = 1'b0; N17 = 1'b1; N21 = 1'b1; N24 = 1'b0; N27 = 1'b0; N30 = 1'b0; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b1; N47 = 1'b1; N50 = 1'b1; N53 = 1'b1; N56 = 1'b0; N60 = 1'b0; N63 = 1'b1; N66 = 1'b1; N69 = 1'b1; N73 = 1'b0; N76 = 1'b1; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b1; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b1; N108 = 1'b1; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b1; N11 = 1'b1; N14 = 1'b1; N17 = 1'b1; N21 = 1'b1; N24 = 1'b1; N27 = 1'b1; N30 = 1'b0; N34 = 1'b1; N37 = 1'b1; N40 = 1'b1; N43 = 1'b1; N47 = 1'b1; N50 = 1'b0; N53 = 1'b1; N56 = 1'b0; N60 = 1'b0; N63 = 1'b1; N66 = 1'b1; N69 = 1'b0; N73 = 1'b1; N76 = 1'b0; N79 = 1'b0; N82 = 1'b0; N86 = 1'b0; N89 = 1'b0; N92 = 1'b0; N95 = 1'b1; N99 = 1'b1; N102 = 1'b1; N105 = 1'b0; N108 = 1'b0; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b0; N8 = 1'b0; N11 = 1'b0; N14 = 1'b0; N17 = 1'b0; N21 = 1'b0; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b1; N37 = 1'b1; N40 = 1'b0; N43 = 1'b1; N47 = 1'b1; N50 = 1'b0; N53 = 1'b1; N56 = 1'b1; N60 = 1'b1; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b0; N76 = 1'b1; N79 = 1'b1; N82 = 1'b0; N86 = 1'b1; N89 = 1'b0; N92 = 1'b1; N95 = 1'b1; N99 = 1'b1; N102 = 1'b1; N105 = 1'b1; N108 = 1'b1; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b0; N8 = 1'b1; N11 = 1'b0; N14 = 1'b0; N17 = 1'b1; N21 = 1'b1; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b0; N37 = 1'b1; N40 = 1'b1; N43 = 1'b1; N47 = 1'b1; N50 = 1'b1; N53 = 1'b0; N56 = 1'b1; N60 = 1'b1; N63 = 1'b1; N66 = 1'b0; N69 = 1'b0; N73 = 1'b0; N76 = 1'b1; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b1; N92 = 1'b1; N95 = 1'b0; N99 = 1'b0; N102 = 1'b0; N105 = 1'b0; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b1; N11 = 1'b0; N14 = 1'b1; N17 = 1'b0; N21 = 1'b0; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b0; N37 = 1'b1; N40 = 1'b1; N43 = 1'b0; N47 = 1'b1; N50 = 1'b1; N53 = 1'b0; N56 = 1'b0; N60 = 1'b0; N63 = 1'b0; N66 = 1'b1; N69 = 1'b1; N73 = 1'b0; N76 = 1'b1; N79 = 1'b1; N82 = 1'b0; N86 = 1'b1; N89 = 1'b1; N92 = 1'b0; N95 = 1'b0; N99 = 1'b1; N102 = 1'b1; N105 = 1'b1; N108 = 1'b0; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b0; N8 = 1'b0; N11 = 1'b1; N14 = 1'b0; N17 = 1'b0; N21 = 1'b0; N24 = 1'b1; N27 = 1'b1; N30 = 1'b0; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b1; N47 = 1'b0; N50 = 1'b0; N53 = 1'b1; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b1; N69 = 1'b1; N73 = 1'b1; N76 = 1'b1; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b1; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b1; N105 = 1'b1; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b0; N11 = 1'b1; N14 = 1'b1; N17 = 1'b0; N21 = 1'b1; N24 = 1'b0; N27 = 1'b0; N30 = 1'b0; N34 = 1'b1; N37 = 1'b0; N40 = 1'b1; N43 = 1'b0; N47 = 1'b0; N50 = 1'b1; N53 = 1'b0; N56 = 1'b1; N60 = 1'b1; N63 = 1'b0; N66 = 1'b1; N69 = 1'b1; N73 = 1'b1; N76 = 1'b1; N79 = 1'b0; N82 = 1'b0; N86 = 1'b0; N89 = 1'b0; N92 = 1'b0; N95 = 1'b0; N99 = 1'b0; N102 = 1'b1; N105 = 1'b0; N108 = 1'b1; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b0; N8 = 1'b0; N11 = 1'b0; N14 = 1'b1; N17 = 1'b1; N21 = 1'b1; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b0; N37 = 1'b1; N40 = 1'b0; N43 = 1'b1; N47 = 1'b0; N50 = 1'b0; N53 = 1'b0; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b1; N69 = 1'b1; N73 = 1'b0; N76 = 1'b0; N79 = 1'b0; N82 = 1'b0; N86 = 1'b0; N89 = 1'b1; N92 = 1'b1; N95 = 1'b0; N99 = 1'b0; N102 = 1'b1; N105 = 1'b1; N108 = 1'b0; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b1; N11 = 1'b0; N14 = 1'b0; N17 = 1'b1; N21 = 1'b0; N24 = 1'b1; N27 = 1'b1; N30 = 1'b0; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b0; N47 = 1'b1; N50 = 1'b1; N53 = 1'b0; N56 = 1'b1; N60 = 1'b1; N63 = 1'b0; N66 = 1'b0; N69 = 1'b0; N73 = 1'b1; N76 = 1'b1; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b1; N92 = 1'b1; N95 = 1'b0; N99 = 1'b0; N102 = 1'b1; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b0; N11 = 1'b0; N14 = 1'b1; N17 = 1'b0; N21 = 1'b0; N24 = 1'b1; N27 = 1'b0; N30 = 1'b1; N34 = 1'b0; N37 = 1'b0; N40 = 1'b0; N43 = 1'b0; N47 = 1'b0; N50 = 1'b0; N53 = 1'b1; N56 = 1'b0; N60 = 1'b0; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b0; N76 = 1'b1; N79 = 1'b1; N82 = 1'b0; N86 = 1'b0; N89 = 1'b1; N92 = 1'b0; N95 = 1'b1; N99 = 1'b1; N102 = 1'b1; N105 = 1'b0; N108 = 1'b0; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b1; N11 = 1'b0; N14 = 1'b0; N17 = 1'b1; N21 = 1'b0; N24 = 1'b1; N27 = 1'b1; N30 = 1'b1; N34 = 1'b0; N37 = 1'b0; N40 = 1'b1; N43 = 1'b1; N47 = 1'b0; N50 = 1'b0; N53 = 1'b0; N56 = 1'b0; N60 = 1'b1; N63 = 1'b0; N66 = 1'b1; N69 = 1'b1; N73 = 1'b1; N76 = 1'b0; N79 = 1'b0; N82 = 1'b1; N86 = 1'b0; N89 = 1'b0; N92 = 1'b0; N95 = 1'b1; N99 = 1'b1; N102 = 1'b0; N105 = 1'b1; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b0; N11 = 1'b1; N14 = 1'b0; N17 = 1'b1; N21 = 1'b0; N24 = 1'b0; N27 = 1'b0; N30 = 1'b0; N34 = 1'b0; N37 = 1'b1; N40 = 1'b1; N43 = 1'b0; N47 = 1'b0; N50 = 1'b0; N53 = 1'b1; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b0; N69 = 1'b0; N73 = 1'b1; N76 = 1'b0; N79 = 1'b1; N82 = 1'b0; N86 = 1'b1; N89 = 1'b0; N92 = 1'b0; N95 = 1'b0; N99 = 1'b0; N102 = 1'b0; N105 = 1'b1; N108 = 1'b1; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b1; N11 = 1'b0; N14 = 1'b1; N17 = 1'b0; N21 = 1'b0; N24 = 1'b1; N27 = 1'b0; N30 = 1'b1; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b0; N47 = 1'b1; N50 = 1'b1; N53 = 1'b0; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b1; N69 = 1'b0; N73 = 1'b1; N76 = 1'b0; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b1; N92 = 1'b1; N95 = 1'b0; N99 = 1'b1; N102 = 1'b1; N105 = 1'b1; N108 = 1'b0; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b1; N11 = 1'b1; N14 = 1'b1; N17 = 1'b0; N21 = 1'b0; N24 = 1'b0; N27 = 1'b0; N30 = 1'b0; N34 = 1'b0; N37 = 1'b1; N40 = 1'b1; N43 = 1'b1; N47 = 1'b0; N50 = 1'b1; N53 = 1'b0; N56 = 1'b1; N60 = 1'b0; N63 = 1'b1; N66 = 1'b1; N69 = 1'b1; N73 = 1'b0; N76 = 1'b1; N79 = 1'b0; N82 = 1'b0; N86 = 1'b1; N89 = 1'b1; N92 = 1'b1; N95 = 1'b1; N99 = 1'b0; N102 = 1'b1; N105 = 1'b1; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b0; N11 = 1'b0; N14 = 1'b1; N17 = 1'b1; N21 = 1'b1; N24 = 1'b0; N27 = 1'b0; N30 = 1'b1; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b1; N47 = 1'b1; N50 = 1'b1; N53 = 1'b1; N56 = 1'b1; N60 = 1'b0; N63 = 1'b1; N66 = 1'b0; N69 = 1'b1; N73 = 1'b1; N76 = 1'b0; N79 = 1'b1; N82 = 1'b0; N86 = 1'b1; N89 = 1'b1; N92 = 1'b1; N95 = 1'b0; N99 = 1'b0; N102 = 1'b1; N105 = 1'b0; N108 = 1'b1; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b1; N11 = 1'b1; N14 = 1'b1; N17 = 1'b0; N21 = 1'b0; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b0; N37 = 1'b1; N40 = 1'b0; N43 = 1'b1; N47 = 1'b0; N50 = 1'b1; N53 = 1'b0; N56 = 1'b0; N60 = 1'b1; N63 = 1'b1; N66 = 1'b0; N69 = 1'b1; N73 = 1'b1; N76 = 1'b0; N79 = 1'b1; N82 = 1'b0; N86 = 1'b0; N89 = 1'b1; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b1; N105 = 1'b1; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b1; N11 = 1'b0; N14 = 1'b0; N17 = 1'b0; N21 = 1'b1; N24 = 1'b1; N27 = 1'b0; N30 = 1'b0; N34 = 1'b0; N37 = 1'b0; N40 = 1'b0; N43 = 1'b1; N47 = 1'b1; N50 = 1'b0; N53 = 1'b1; N56 = 1'b1; N60 = 1'b1; N63 = 1'b1; N66 = 1'b0; N69 = 1'b0; N73 = 1'b0; N76 = 1'b1; N79 = 1'b0; N82 = 1'b1; N86 = 1'b1; N89 = 1'b1; N92 = 1'b1; N95 = 1'b1; N99 = 1'b1; N102 = 1'b0; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b1; N11 = 1'b0; N14 = 1'b1; N17 = 1'b1; N21 = 1'b0; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b0; N37 = 1'b1; N40 = 1'b0; N43 = 1'b0; N47 = 1'b0; N50 = 1'b0; N53 = 1'b0; N56 = 1'b1; N60 = 1'b0; N63 = 1'b1; N66 = 1'b0; N69 = 1'b0; N73 = 1'b1; N76 = 1'b1; N79 = 1'b0; N82 = 1'b0; N86 = 1'b1; N89 = 1'b0; N92 = 1'b1; N95 = 1'b1; N99 = 1'b1; N102 = 1'b0; N105 = 1'b0; N108 = 1'b0; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b0; N11 = 1'b1; N14 = 1'b0; N17 = 1'b0; N21 = 1'b0; N24 = 1'b0; N27 = 1'b0; N30 = 1'b1; N34 = 1'b0; N37 = 1'b1; N40 = 1'b0; N43 = 1'b0; N47 = 1'b1; N50 = 1'b1; N53 = 1'b1; N56 = 1'b1; N60 = 1'b0; N63 = 1'b1; N66 = 1'b0; N69 = 1'b0; N73 = 1'b0; N76 = 1'b0; N79 = 1'b0; N82 = 1'b0; N86 = 1'b0; N89 = 1'b1; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b0; N108 = 1'b1; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b1; N11 = 1'b1; N14 = 1'b0; N17 = 1'b0; N21 = 1'b0; N24 = 1'b0; N27 = 1'b1; N30 = 1'b0; N34 = 1'b0; N37 = 1'b1; N40 = 1'b1; N43 = 1'b0; N47 = 1'b1; N50 = 1'b1; N53 = 1'b0; N56 = 1'b0; N60 = 1'b0; N63 = 1'b0; N66 = 1'b0; N69 = 1'b0; N73 = 1'b0; N76 = 1'b1; N79 = 1'b1; N82 = 1'b1; N86 = 1'b1; N89 = 1'b1; N92 = 1'b1; N95 = 1'b0; N99 = 1'b1; N102 = 1'b1; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b0; N11 = 1'b0; N14 = 1'b0; N17 = 1'b0; N21 = 1'b0; N24 = 1'b1; N27 = 1'b0; N30 = 1'b0; N34 = 1'b1; N37 = 1'b1; N40 = 1'b0; N43 = 1'b1; N47 = 1'b1; N50 = 1'b0; N53 = 1'b1; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b1; N69 = 1'b0; N73 = 1'b0; N76 = 1'b0; N79 = 1'b0; N82 = 1'b1; N86 = 1'b1; N89 = 1'b1; N92 = 1'b1; N95 = 1'b0; N99 = 1'b1; N102 = 1'b0; N105 = 1'b0; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b1; N11 = 1'b0; N14 = 1'b1; N17 = 1'b1; N21 = 1'b1; N24 = 1'b1; N27 = 1'b1; N30 = 1'b0; N34 = 1'b1; N37 = 1'b1; N40 = 1'b0; N43 = 1'b1; N47 = 1'b0; N50 = 1'b0; N53 = 1'b0; N56 = 1'b1; N60 = 1'b1; N63 = 1'b1; N66 = 1'b1; N69 = 1'b0; N73 = 1'b1; N76 = 1'b1; N79 = 1'b1; N82 = 1'b0; N86 = 1'b1; N89 = 1'b1; N92 = 1'b0; N95 = 1'b0; N99 = 1'b0; N102 = 1'b0; N105 = 1'b1; N108 = 1'b0; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b0; N11 = 1'b0; N14 = 1'b0; N17 = 1'b0; N21 = 1'b1; N24 = 1'b1; N27 = 1'b0; N30 = 1'b0; N34 = 1'b1; N37 = 1'b0; N40 = 1'b1; N43 = 1'b0; N47 = 1'b1; N50 = 1'b1; N53 = 1'b1; N56 = 1'b0; N60 = 1'b1; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b1; N76 = 1'b0; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b1; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b1; N105 = 1'b1; N108 = 1'b0; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b0; N11 = 1'b1; N14 = 1'b0; N17 = 1'b1; N21 = 1'b0; N24 = 1'b0; N27 = 1'b0; N30 = 1'b1; N34 = 1'b1; N37 = 1'b0; N40 = 1'b1; N43 = 1'b0; N47 = 1'b0; N50 = 1'b1; N53 = 1'b0; N56 = 1'b0; N60 = 1'b0; N63 = 1'b1; N66 = 1'b1; N69 = 1'b0; N73 = 1'b1; N76 = 1'b1; N79 = 1'b1; N82 = 1'b0; N86 = 1'b0; N89 = 1'b1; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b1; N105 = 1'b0; N108 = 1'b0; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b1; N11 = 1'b0; N14 = 1'b0; N17 = 1'b0; N21 = 1'b1; N24 = 1'b0; N27 = 1'b1; N30 = 1'b0; N34 = 1'b0; N37 = 1'b1; N40 = 1'b1; N43 = 1'b0; N47 = 1'b0; N50 = 1'b0; N53 = 1'b0; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b1; N69 = 1'b0; N73 = 1'b1; N76 = 1'b0; N79 = 1'b0; N82 = 1'b0; N86 = 1'b1; N89 = 1'b1; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b1; N11 = 1'b1; N14 = 1'b0; N17 = 1'b0; N21 = 1'b1; N24 = 1'b0; N27 = 1'b0; N30 = 1'b1; N34 = 1'b0; N37 = 1'b1; N40 = 1'b1; N43 = 1'b1; N47 = 1'b1; N50 = 1'b1; N53 = 1'b1; N56 = 1'b1; N60 = 1'b1; N63 = 1'b1; N66 = 1'b0; N69 = 1'b0; N73 = 1'b1; N76 = 1'b0; N79 = 1'b1; N82 = 1'b1; N86 = 1'b1; N89 = 1'b0; N92 = 1'b1; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b1; N108 = 1'b0; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b1; N11 = 1'b0; N14 = 1'b0; N17 = 1'b0; N21 = 1'b1; N24 = 1'b0; N27 = 1'b0; N30 = 1'b0; N34 = 1'b1; N37 = 1'b1; N40 = 1'b0; N43 = 1'b1; N47 = 1'b1; N50 = 1'b0; N53 = 1'b0; N56 = 1'b1; N60 = 1'b1; N63 = 1'b1; N66 = 1'b1; N69 = 1'b1; N73 = 1'b1; N76 = 1'b0; N79 = 1'b0; N82 = 1'b0; N86 = 1'b1; N89 = 1'b1; N92 = 1'b0; N95 = 1'b0; N99 = 1'b0; N102 = 1'b1; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b0; N11 = 1'b1; N14 = 1'b0; N17 = 1'b1; N21 = 1'b0; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b0; N37 = 1'b0; N40 = 1'b0; N43 = 1'b0; N47 = 1'b0; N50 = 1'b0; N53 = 1'b1; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b1; N76 = 1'b0; N79 = 1'b0; N82 = 1'b0; N86 = 1'b1; N89 = 1'b1; N92 = 1'b1; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b0; N108 = 1'b0; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b0; N11 = 1'b0; N14 = 1'b0; N17 = 1'b1; N21 = 1'b1; N24 = 1'b1; N27 = 1'b0; N30 = 1'b1; N34 = 1'b0; N37 = 1'b0; N40 = 1'b0; N43 = 1'b0; N47 = 1'b0; N50 = 1'b0; N53 = 1'b0; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b0; N69 = 1'b0; N73 = 1'b1; N76 = 1'b1; N79 = 1'b1; N82 = 1'b0; N86 = 1'b1; N89 = 1'b1; N92 = 1'b1; N95 = 1'b0; N99 = 1'b1; N102 = 1'b0; N105 = 1'b1; N108 = 1'b0; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b0; N11 = 1'b1; N14 = 1'b0; N17 = 1'b1; N21 = 1'b0; N24 = 1'b1; N27 = 1'b0; N30 = 1'b1; N34 = 1'b1; N37 = 1'b1; N40 = 1'b1; N43 = 1'b0; N47 = 1'b1; N50 = 1'b1; N53 = 1'b1; N56 = 1'b0; N60 = 1'b1; N63 = 1'b0; N66 = 1'b0; N69 = 1'b0; N73 = 1'b0; N76 = 1'b1; N79 = 1'b1; N82 = 1'b0; N86 = 1'b1; N89 = 1'b1; N92 = 1'b1; N95 = 1'b0; N99 = 1'b0; N102 = 1'b1; N105 = 1'b0; N108 = 1'b0; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b0; N11 = 1'b1; N14 = 1'b1; N17 = 1'b0; N21 = 1'b1; N24 = 1'b1; N27 = 1'b0; N30 = 1'b0; N34 = 1'b1; N37 = 1'b0; N40 = 1'b1; N43 = 1'b0; N47 = 1'b0; N50 = 1'b1; N53 = 1'b1; N56 = 1'b1; N60 = 1'b0; N63 = 1'b1; N66 = 1'b0; N69 = 1'b0; N73 = 1'b0; N76 = 1'b1; N79 = 1'b0; N82 = 1'b1; N86 = 1'b0; N89 = 1'b1; N92 = 1'b0; N95 = 1'b1; N99 = 1'b1; N102 = 1'b0; N105 = 1'b1; N108 = 1'b0; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b0; N11 = 1'b0; N14 = 1'b1; N17 = 1'b0; N21 = 1'b0; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b0; N37 = 1'b0; N40 = 1'b0; N43 = 1'b1; N47 = 1'b1; N50 = 1'b0; N53 = 1'b1; N56 = 1'b0; N60 = 1'b1; N63 = 1'b1; N66 = 1'b0; N69 = 1'b0; N73 = 1'b1; N76 = 1'b0; N79 = 1'b0; N82 = 1'b1; N86 = 1'b0; N89 = 1'b1; N92 = 1'b1; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b1; N108 = 1'b1; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b0; N11 = 1'b0; N14 = 1'b1; N17 = 1'b1; N21 = 1'b1; N24 = 1'b1; N27 = 1'b0; N30 = 1'b0; N34 = 1'b1; N37 = 1'b1; N40 = 1'b0; N43 = 1'b0; N47 = 1'b0; N50 = 1'b1; N53 = 1'b1; N56 = 1'b0; N60 = 1'b0; N63 = 1'b0; N66 = 1'b0; N69 = 1'b0; N73 = 1'b1; N76 = 1'b0; N79 = 1'b0; N82 = 1'b0; N86 = 1'b0; N89 = 1'b1; N92 = 1'b1; N95 = 1'b1; N99 = 1'b1; N102 = 1'b1; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b1; N11 = 1'b0; N14 = 1'b1; N17 = 1'b1; N21 = 1'b0; N24 = 1'b1; N27 = 1'b0; N30 = 1'b1; N34 = 1'b1; N37 = 1'b1; N40 = 1'b1; N43 = 1'b1; N47 = 1'b1; N50 = 1'b1; N53 = 1'b0; N56 = 1'b1; N60 = 1'b1; N63 = 1'b1; N66 = 1'b1; N69 = 1'b1; N73 = 1'b1; N76 = 1'b1; N79 = 1'b1; N82 = 1'b0; N86 = 1'b1; N89 = 1'b1; N92 = 1'b0; N95 = 1'b0; N99 = 1'b0; N102 = 1'b1; N105 = 1'b1; N108 = 1'b0; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b0; N11 = 1'b0; N14 = 1'b1; N17 = 1'b0; N21 = 1'b0; N24 = 1'b0; N27 = 1'b0; N30 = 1'b0; N34 = 1'b0; N37 = 1'b1; N40 = 1'b1; N43 = 1'b0; N47 = 1'b1; N50 = 1'b1; N53 = 1'b0; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b1; N69 = 1'b1; N73 = 1'b1; N76 = 1'b1; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b0; N92 = 1'b0; N95 = 1'b0; N99 = 1'b0; N102 = 1'b0; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b0; N11 = 1'b1; N14 = 1'b0; N17 = 1'b1; N21 = 1'b1; N24 = 1'b1; N27 = 1'b1; N30 = 1'b1; N34 = 1'b0; N37 = 1'b1; N40 = 1'b0; N43 = 1'b1; N47 = 1'b0; N50 = 1'b0; N53 = 1'b0; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b0; N76 = 1'b0; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b0; N92 = 1'b1; N95 = 1'b1; N99 = 1'b0; N102 = 1'b1; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b0; N8 = 1'b0; N11 = 1'b0; N14 = 1'b1; N17 = 1'b1; N21 = 1'b0; N24 = 1'b0; N27 = 1'b0; N30 = 1'b0; N34 = 1'b1; N37 = 1'b1; N40 = 1'b0; N43 = 1'b1; N47 = 1'b1; N50 = 1'b1; N53 = 1'b0; N56 = 1'b1; N60 = 1'b1; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b0; N76 = 1'b0; N79 = 1'b0; N82 = 1'b1; N86 = 1'b1; N89 = 1'b0; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b1; N105 = 1'b1; N108 = 1'b1; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b0; N8 = 1'b0; N11 = 1'b0; N14 = 1'b1; N17 = 1'b1; N21 = 1'b1; N24 = 1'b0; N27 = 1'b1; N30 = 1'b0; N34 = 1'b1; N37 = 1'b1; N40 = 1'b1; N43 = 1'b1; N47 = 1'b1; N50 = 1'b1; N53 = 1'b1; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b1; N76 = 1'b0; N79 = 1'b0; N82 = 1'b1; N86 = 1'b1; N89 = 1'b0; N92 = 1'b0; N95 = 1'b1; N99 = 1'b1; N102 = 1'b0; N105 = 1'b0; N108 = 1'b0; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b1; N11 = 1'b1; N14 = 1'b0; N17 = 1'b0; N21 = 1'b0; N24 = 1'b0; N27 = 1'b1; N30 = 1'b0; N34 = 1'b1; N37 = 1'b1; N40 = 1'b0; N43 = 1'b0; N47 = 1'b0; N50 = 1'b1; N53 = 1'b1; N56 = 1'b1; N60 = 1'b1; N63 = 1'b1; N66 = 1'b1; N69 = 1'b1; N73 = 1'b0; N76 = 1'b0; N79 = 1'b0; N82 = 1'b1; N86 = 1'b0; N89 = 1'b1; N92 = 1'b1; N95 = 1'b0; N99 = 1'b0; N102 = 1'b1; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b0; N8 = 1'b1; N11 = 1'b1; N14 = 1'b1; N17 = 1'b0; N21 = 1'b0; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b1; N37 = 1'b1; N40 = 1'b1; N43 = 1'b0; N47 = 1'b1; N50 = 1'b0; N53 = 1'b0; N56 = 1'b1; N60 = 1'b0; N63 = 1'b1; N66 = 1'b0; N69 = 1'b1; N73 = 1'b1; N76 = 1'b0; N79 = 1'b1; N82 = 1'b1; N86 = 1'b1; N89 = 1'b1; N92 = 1'b0; N95 = 1'b0; N99 = 1'b1; N102 = 1'b1; N105 = 1'b1; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b1; N11 = 1'b0; N14 = 1'b1; N17 = 1'b0; N21 = 1'b1; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b1; N37 = 1'b0; N40 = 1'b1; N43 = 1'b0; N47 = 1'b0; N50 = 1'b0; N53 = 1'b1; N56 = 1'b1; N60 = 1'b1; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b0; N76 = 1'b1; N79 = 1'b0; N82 = 1'b1; N86 = 1'b1; N89 = 1'b0; N92 = 1'b1; N95 = 1'b0; N99 = 1'b1; N102 = 1'b0; N105 = 1'b0; N108 = 1'b0; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b1; N11 = 1'b0; N14 = 1'b1; N17 = 1'b0; N21 = 1'b1; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b1; N37 = 1'b1; N40 = 1'b0; N43 = 1'b0; N47 = 1'b0; N50 = 1'b0; N53 = 1'b1; N56 = 1'b0; N60 = 1'b0; N63 = 1'b1; N66 = 1'b0; N69 = 1'b1; N73 = 1'b1; N76 = 1'b1; N79 = 1'b0; N82 = 1'b1; N86 = 1'b1; N89 = 1'b0; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b1; N108 = 1'b0; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b0; N8 = 1'b0; N11 = 1'b1; N14 = 1'b1; N17 = 1'b0; N21 = 1'b1; N24 = 1'b0; N27 = 1'b1; N30 = 1'b0; N34 = 1'b0; N37 = 1'b0; N40 = 1'b0; N43 = 1'b1; N47 = 1'b1; N50 = 1'b1; N53 = 1'b0; N56 = 1'b0; N60 = 1'b0; N63 = 1'b1; N66 = 1'b0; N69 = 1'b1; N73 = 1'b1; N76 = 1'b0; N79 = 1'b0; N82 = 1'b1; N86 = 1'b0; N89 = 1'b0; N92 = 1'b1; N95 = 1'b0; N99 = 1'b0; N102 = 1'b0; N105 = 1'b0; N108 = 1'b0; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b0; N11 = 1'b0; N14 = 1'b0; N17 = 1'b1; N21 = 1'b0; N24 = 1'b0; N27 = 1'b0; N30 = 1'b1; N34 = 1'b0; N37 = 1'b1; N40 = 1'b1; N43 = 1'b1; N47 = 1'b1; N50 = 1'b1; N53 = 1'b0; N56 = 1'b0; N60 = 1'b1; N63 = 1'b1; N66 = 1'b1; N69 = 1'b1; N73 = 1'b0; N76 = 1'b1; N79 = 1'b0; N82 = 1'b0; N86 = 1'b1; N89 = 1'b1; N92 = 1'b1; N95 = 1'b0; N99 = 1'b1; N102 = 1'b1; N105 = 1'b0; N108 = 1'b1; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b0; N8 = 1'b1; N11 = 1'b0; N14 = 1'b1; N17 = 1'b0; N21 = 1'b1; N24 = 1'b0; N27 = 1'b0; N30 = 1'b1; N34 = 1'b0; N37 = 1'b0; N40 = 1'b1; N43 = 1'b0; N47 = 1'b0; N50 = 1'b1; N53 = 1'b0; N56 = 1'b0; N60 = 1'b1; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b0; N76 = 1'b1; N79 = 1'b1; N82 = 1'b1; N86 = 1'b1; N89 = 1'b1; N92 = 1'b1; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b1; N108 = 1'b0; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b0; N8 = 1'b1; N11 = 1'b0; N14 = 1'b0; N17 = 1'b1; N21 = 1'b1; N24 = 1'b1; N27 = 1'b0; N30 = 1'b1; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b1; N47 = 1'b1; N50 = 1'b1; N53 = 1'b1; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b1; N69 = 1'b1; N73 = 1'b1; N76 = 1'b1; N79 = 1'b0; N82 = 1'b0; N86 = 1'b1; N89 = 1'b1; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b1; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b0; N11 = 1'b1; N14 = 1'b0; N17 = 1'b0; N21 = 1'b0; N24 = 1'b1; N27 = 1'b0; N30 = 1'b0; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b1; N47 = 1'b0; N50 = 1'b0; N53 = 1'b1; N56 = 1'b0; N60 = 1'b0; N63 = 1'b1; N66 = 1'b1; N69 = 1'b0; N73 = 1'b1; N76 = 1'b1; N79 = 1'b0; N82 = 1'b1; N86 = 1'b1; N89 = 1'b1; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b0; N11 = 1'b0; N14 = 1'b0; N17 = 1'b1; N21 = 1'b1; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b0; N47 = 1'b1; N50 = 1'b0; N53 = 1'b1; N56 = 1'b0; N60 = 1'b0; N63 = 1'b0; N66 = 1'b1; N69 = 1'b1; N73 = 1'b1; N76 = 1'b1; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b1; N92 = 1'b1; N95 = 1'b1; N99 = 1'b1; N102 = 1'b1; N105 = 1'b1; N108 = 1'b0; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b1; N11 = 1'b0; N14 = 1'b0; N17 = 1'b1; N21 = 1'b0; N24 = 1'b1; N27 = 1'b0; N30 = 1'b0; N34 = 1'b0; N37 = 1'b0; N40 = 1'b0; N43 = 1'b1; N47 = 1'b0; N50 = 1'b1; N53 = 1'b1; N56 = 1'b1; N60 = 1'b1; N63 = 1'b1; N66 = 1'b1; N69 = 1'b0; N73 = 1'b1; N76 = 1'b0; N79 = 1'b0; N82 = 1'b1; N86 = 1'b0; N89 = 1'b0; N92 = 1'b0; N95 = 1'b0; N99 = 1'b0; N102 = 1'b1; N105 = 1'b1; N108 = 1'b1; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b0; N11 = 1'b1; N14 = 1'b0; N17 = 1'b1; N21 = 1'b1; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b0; N37 = 1'b0; N40 = 1'b1; N43 = 1'b1; N47 = 1'b0; N50 = 1'b0; N53 = 1'b0; N56 = 1'b0; N60 = 1'b0; N63 = 1'b1; N66 = 1'b1; N69 = 1'b0; N73 = 1'b0; N76 = 1'b0; N79 = 1'b0; N82 = 1'b1; N86 = 1'b0; N89 = 1'b1; N92 = 1'b1; N95 = 1'b0; N99 = 1'b1; N102 = 1'b0; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b0; N11 = 1'b1; N14 = 1'b1; N17 = 1'b1; N21 = 1'b0; N24 = 1'b1; N27 = 1'b1; N30 = 1'b1; N34 = 1'b0; N37 = 1'b1; N40 = 1'b0; N43 = 1'b0; N47 = 1'b0; N50 = 1'b0; N53 = 1'b0; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b1; N69 = 1'b1; N73 = 1'b0; N76 = 1'b1; N79 = 1'b0; N82 = 1'b1; N86 = 1'b0; N89 = 1'b0; N92 = 1'b1; N95 = 1'b0; N99 = 1'b0; N102 = 1'b1; N105 = 1'b0; N108 = 1'b0; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b1; N11 = 1'b0; N14 = 1'b1; N17 = 1'b0; N21 = 1'b1; N24 = 1'b1; N27 = 1'b0; N30 = 1'b1; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b1; N47 = 1'b0; N50 = 1'b0; N53 = 1'b1; N56 = 1'b1; N60 = 1'b1; N63 = 1'b1; N66 = 1'b0; N69 = 1'b1; N73 = 1'b1; N76 = 1'b0; N79 = 1'b0; N82 = 1'b1; N86 = 1'b1; N89 = 1'b0; N92 = 1'b0; N95 = 1'b0; N99 = 1'b0; N102 = 1'b1; N105 = 1'b1; N108 = 1'b0; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b1; N11 = 1'b1; N14 = 1'b1; N17 = 1'b1; N21 = 1'b0; N24 = 1'b1; N27 = 1'b1; N30 = 1'b0; N34 = 1'b0; N37 = 1'b1; N40 = 1'b0; N43 = 1'b0; N47 = 1'b1; N50 = 1'b0; N53 = 1'b0; N56 = 1'b0; N60 = 1'b1; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b0; N76 = 1'b1; N79 = 1'b0; N82 = 1'b0; N86 = 1'b1; N89 = 1'b0; N92 = 1'b0; N95 = 1'b0; N99 = 1'b1; N102 = 1'b0; N105 = 1'b0; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b0; N11 = 1'b0; N14 = 1'b1; N17 = 1'b0; N21 = 1'b0; N24 = 1'b1; N27 = 1'b0; N30 = 1'b0; N34 = 1'b0; N37 = 1'b0; N40 = 1'b1; N43 = 1'b0; N47 = 1'b1; N50 = 1'b0; N53 = 1'b0; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b0; N76 = 1'b1; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b0; N92 = 1'b1; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b0; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b0; N8 = 1'b1; N11 = 1'b1; N14 = 1'b1; N17 = 1'b1; N21 = 1'b1; N24 = 1'b1; N27 = 1'b1; N30 = 1'b1; N34 = 1'b0; N37 = 1'b1; N40 = 1'b0; N43 = 1'b0; N47 = 1'b0; N50 = 1'b1; N53 = 1'b1; N56 = 1'b1; N60 = 1'b1; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b0; N76 = 1'b1; N79 = 1'b0; N82 = 1'b1; N86 = 1'b0; N89 = 1'b1; N92 = 1'b0; N95 = 1'b1; N99 = 1'b1; N102 = 1'b1; N105 = 1'b1; N108 = 1'b0; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b1; N11 = 1'b1; N14 = 1'b1; N17 = 1'b1; N21 = 1'b1; N24 = 1'b0; N27 = 1'b0; N30 = 1'b1; N34 = 1'b0; N37 = 1'b0; N40 = 1'b0; N43 = 1'b0; N47 = 1'b1; N50 = 1'b1; N53 = 1'b1; N56 = 1'b0; N60 = 1'b1; N63 = 1'b0; N66 = 1'b1; N69 = 1'b1; N73 = 1'b1; N76 = 1'b0; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b1; N92 = 1'b0; N95 = 1'b0; N99 = 1'b0; N102 = 1'b1; N105 = 1'b1; N108 = 1'b1; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b1; N11 = 1'b0; N14 = 1'b0; N17 = 1'b1; N21 = 1'b1; N24 = 1'b1; N27 = 1'b0; N30 = 1'b1; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b1; N47 = 1'b1; N50 = 1'b1; N53 = 1'b0; N56 = 1'b0; N60 = 1'b1; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b1; N76 = 1'b1; N79 = 1'b0; N82 = 1'b1; N86 = 1'b1; N89 = 1'b0; N92 = 1'b0; N95 = 1'b0; N99 = 1'b0; N102 = 1'b0; N105 = 1'b1; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b1; N11 = 1'b1; N14 = 1'b0; N17 = 1'b1; N21 = 1'b0; N24 = 1'b0; N27 = 1'b1; N30 = 1'b0; N34 = 1'b0; N37 = 1'b0; N40 = 1'b0; N43 = 1'b0; N47 = 1'b0; N50 = 1'b1; N53 = 1'b1; N56 = 1'b0; N60 = 1'b1; N63 = 1'b1; N66 = 1'b1; N69 = 1'b0; N73 = 1'b0; N76 = 1'b0; N79 = 1'b0; N82 = 1'b1; N86 = 1'b0; N89 = 1'b0; N92 = 1'b1; N95 = 1'b1; N99 = 1'b1; N102 = 1'b1; N105 = 1'b0; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b0; N11 = 1'b1; N14 = 1'b0; N17 = 1'b0; N21 = 1'b1; N24 = 1'b0; N27 = 1'b0; N30 = 1'b1; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b0; N47 = 1'b1; N50 = 1'b0; N53 = 1'b0; N56 = 1'b1; N60 = 1'b0; N63 = 1'b1; N66 = 1'b0; N69 = 1'b0; N73 = 1'b1; N76 = 1'b1; N79 = 1'b0; N82 = 1'b1; N86 = 1'b1; N89 = 1'b1; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b0; N11 = 1'b1; N14 = 1'b1; N17 = 1'b0; N21 = 1'b1; N24 = 1'b0; N27 = 1'b1; N30 = 1'b0; N34 = 1'b1; N37 = 1'b1; N40 = 1'b1; N43 = 1'b0; N47 = 1'b1; N50 = 1'b0; N53 = 1'b0; N56 = 1'b0; N60 = 1'b1; N63 = 1'b1; N66 = 1'b1; N69 = 1'b1; N73 = 1'b0; N76 = 1'b1; N79 = 1'b1; N82 = 1'b0; N86 = 1'b1; N89 = 1'b0; N92 = 1'b1; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b1; N108 = 1'b1; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b0; N11 = 1'b0; N14 = 1'b0; N17 = 1'b0; N21 = 1'b0; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b0; N37 = 1'b0; N40 = 1'b1; N43 = 1'b0; N47 = 1'b0; N50 = 1'b0; N53 = 1'b0; N56 = 1'b0; N60 = 1'b1; N63 = 1'b1; N66 = 1'b0; N69 = 1'b1; N73 = 1'b1; N76 = 1'b1; N79 = 1'b0; N82 = 1'b0; N86 = 1'b1; N89 = 1'b0; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b1; N105 = 1'b1; N108 = 1'b0; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b0; N11 = 1'b1; N14 = 1'b1; N17 = 1'b0; N21 = 1'b0; N24 = 1'b1; N27 = 1'b0; N30 = 1'b1; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b1; N47 = 1'b0; N50 = 1'b1; N53 = 1'b1; N56 = 1'b0; N60 = 1'b1; N63 = 1'b0; N66 = 1'b1; N69 = 1'b1; N73 = 1'b1; N76 = 1'b0; N79 = 1'b1; N82 = 1'b0; N86 = 1'b0; N89 = 1'b0; N92 = 1'b1; N95 = 1'b0; N99 = 1'b1; N102 = 1'b1; N105 = 1'b1; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b0; N11 = 1'b0; N14 = 1'b0; N17 = 1'b1; N21 = 1'b0; N24 = 1'b1; N27 = 1'b1; N30 = 1'b1; N34 = 1'b1; N37 = 1'b0; N40 = 1'b1; N43 = 1'b1; N47 = 1'b1; N50 = 1'b0; N53 = 1'b0; N56 = 1'b1; N60 = 1'b1; N63 = 1'b0; N66 = 1'b0; N69 = 1'b0; N73 = 1'b1; N76 = 1'b0; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b0; N92 = 1'b1; N95 = 1'b1; N99 = 1'b0; N102 = 1'b1; N105 = 1'b0; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b0; N11 = 1'b0; N14 = 1'b0; N17 = 1'b0; N21 = 1'b1; N24 = 1'b0; N27 = 1'b1; N30 = 1'b0; N34 = 1'b0; N37 = 1'b0; N40 = 1'b0; N43 = 1'b1; N47 = 1'b1; N50 = 1'b0; N53 = 1'b0; N56 = 1'b0; N60 = 1'b0; N63 = 1'b0; N66 = 1'b1; N69 = 1'b1; N73 = 1'b1; N76 = 1'b1; N79 = 1'b1; N82 = 1'b0; N86 = 1'b0; N89 = 1'b0; N92 = 1'b1; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b0; N108 = 1'b1; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b1; N11 = 1'b1; N14 = 1'b0; N17 = 1'b0; N21 = 1'b0; N24 = 1'b1; N27 = 1'b1; N30 = 1'b0; N34 = 1'b1; N37 = 1'b0; N40 = 1'b1; N43 = 1'b1; N47 = 1'b1; N50 = 1'b0; N53 = 1'b1; N56 = 1'b1; N60 = 1'b0; N63 = 1'b1; N66 = 1'b0; N69 = 1'b0; N73 = 1'b1; N76 = 1'b0; N79 = 1'b1; N82 = 1'b1; N86 = 1'b1; N89 = 1'b0; N92 = 1'b0; N95 = 1'b1; N99 = 1'b1; N102 = 1'b1; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b1; N11 = 1'b0; N14 = 1'b1; N17 = 1'b1; N21 = 1'b1; N24 = 1'b0; N27 = 1'b0; N30 = 1'b1; N34 = 1'b0; N37 = 1'b0; N40 = 1'b1; N43 = 1'b0; N47 = 1'b0; N50 = 1'b1; N53 = 1'b0; N56 = 1'b1; N60 = 1'b1; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b1; N76 = 1'b0; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b1; N92 = 1'b0; N95 = 1'b0; N99 = 1'b0; N102 = 1'b0; N105 = 1'b1; N108 = 1'b1; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b0; N11 = 1'b1; N14 = 1'b1; N17 = 1'b0; N21 = 1'b0; N24 = 1'b1; N27 = 1'b0; N30 = 1'b1; N34 = 1'b0; N37 = 1'b0; N40 = 1'b1; N43 = 1'b1; N47 = 1'b0; N50 = 1'b1; N53 = 1'b0; N56 = 1'b1; N60 = 1'b1; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b0; N76 = 1'b1; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b1; N92 = 1'b1; N95 = 1'b1; N99 = 1'b1; N102 = 1'b0; N105 = 1'b1; N108 = 1'b1; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b1; N11 = 1'b1; N14 = 1'b0; N17 = 1'b1; N21 = 1'b0; N24 = 1'b0; N27 = 1'b0; N30 = 1'b1; N34 = 1'b0; N37 = 1'b0; N40 = 1'b1; N43 = 1'b1; N47 = 1'b1; N50 = 1'b0; N53 = 1'b1; N56 = 1'b0; N60 = 1'b0; N63 = 1'b0; N66 = 1'b0; N69 = 1'b0; N73 = 1'b0; N76 = 1'b0; N79 = 1'b1; N82 = 1'b0; N86 = 1'b0; N89 = 1'b0; N92 = 1'b0; N95 = 1'b0; N99 = 1'b0; N102 = 1'b1; N105 = 1'b0; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b0; N8 = 1'b1; N11 = 1'b1; N14 = 1'b1; N17 = 1'b0; N21 = 1'b1; N24 = 1'b1; N27 = 1'b1; N30 = 1'b0; N34 = 1'b0; N37 = 1'b1; N40 = 1'b0; N43 = 1'b1; N47 = 1'b1; N50 = 1'b0; N53 = 1'b0; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b0; N69 = 1'b0; N73 = 1'b0; N76 = 1'b0; N79 = 1'b1; N82 = 1'b0; N86 = 1'b0; N89 = 1'b1; N92 = 1'b0; N95 = 1'b0; N99 = 1'b1; N102 = 1'b0; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b0; N11 = 1'b1; N14 = 1'b0; N17 = 1'b1; N21 = 1'b0; N24 = 1'b1; N27 = 1'b1; N30 = 1'b1; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b1; N47 = 1'b0; N50 = 1'b0; N53 = 1'b0; N56 = 1'b0; N60 = 1'b0; N63 = 1'b1; N66 = 1'b0; N69 = 1'b1; N73 = 1'b0; N76 = 1'b0; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b1; N92 = 1'b1; N95 = 1'b0; N99 = 1'b0; N102 = 1'b0; N105 = 1'b0; N108 = 1'b1; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b1; N11 = 1'b0; N14 = 1'b0; N17 = 1'b0; N21 = 1'b0; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b0; N47 = 1'b0; N50 = 1'b0; N53 = 1'b1; N56 = 1'b0; N60 = 1'b1; N63 = 1'b1; N66 = 1'b0; N69 = 1'b0; N73 = 1'b0; N76 = 1'b1; N79 = 1'b0; N82 = 1'b0; N86 = 1'b1; N89 = 1'b1; N92 = 1'b0; N95 = 1'b0; N99 = 1'b0; N102 = 1'b1; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b0; N11 = 1'b0; N14 = 1'b1; N17 = 1'b0; N21 = 1'b0; N24 = 1'b0; N27 = 1'b1; N30 = 1'b1; N34 = 1'b1; N37 = 1'b1; N40 = 1'b1; N43 = 1'b0; N47 = 1'b1; N50 = 1'b0; N53 = 1'b1; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b1; N76 = 1'b0; N79 = 1'b1; N82 = 1'b1; N86 = 1'b1; N89 = 1'b1; N92 = 1'b0; N95 = 1'b0; N99 = 1'b0; N102 = 1'b1; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b1; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b0; N11 = 1'b1; N14 = 1'b0; N17 = 1'b1; N21 = 1'b1; N24 = 1'b0; N27 = 1'b1; N30 = 1'b0; N34 = 1'b1; N37 = 1'b1; N40 = 1'b0; N43 = 1'b1; N47 = 1'b1; N50 = 1'b1; N53 = 1'b1; N56 = 1'b1; N60 = 1'b0; N63 = 1'b0; N66 = 1'b1; N69 = 1'b0; N73 = 1'b1; N76 = 1'b1; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b0; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b1; N105 = 1'b0; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b0; N11 = 1'b0; N14 = 1'b1; N17 = 1'b1; N21 = 1'b1; N24 = 1'b0; N27 = 1'b0; N30 = 1'b1; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b1; N47 = 1'b1; N50 = 1'b0; N53 = 1'b0; N56 = 1'b0; N60 = 1'b0; N63 = 1'b0; N66 = 1'b0; N69 = 1'b0; N73 = 1'b1; N76 = 1'b1; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b0; N92 = 1'b1; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b1; N108 = 1'b1; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b1; N11 = 1'b1; N14 = 1'b0; N17 = 1'b0; N21 = 1'b0; N24 = 1'b1; N27 = 1'b1; N30 = 1'b0; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b0; N47 = 1'b0; N50 = 1'b1; N53 = 1'b0; N56 = 1'b1; N60 = 1'b0; N63 = 1'b1; N66 = 1'b0; N69 = 1'b1; N73 = 1'b0; N76 = 1'b0; N79 = 1'b1; N82 = 1'b0; N86 = 1'b1; N89 = 1'b1; N92 = 1'b0; N95 = 1'b1; N99 = 1'b0; N102 = 1'b0; N105 = 1'b1; N108 = 1'b0; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b0; N11 = 1'b1; N14 = 1'b1; N17 = 1'b0; N21 = 1'b0; N24 = 1'b1; N27 = 1'b0; N30 = 1'b0; N34 = 1'b1; N37 = 1'b1; N40 = 1'b0; N43 = 1'b1; N47 = 1'b1; N50 = 1'b0; N53 = 1'b0; N56 = 1'b1; N60 = 1'b1; N63 = 1'b0; N66 = 1'b0; N69 = 1'b1; N73 = 1'b0; N76 = 1'b1; N79 = 1'b0; N82 = 1'b0; N86 = 1'b1; N89 = 1'b1; N92 = 1'b1; N95 = 1'b1; N99 = 1'b0; N102 = 1'b1; N105 = 1'b1; N108 = 1'b0; N112 = 1'b0; N115 = 1'b1; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b0; N11 = 1'b0; N14 = 1'b0; N17 = 1'b1; N21 = 1'b1; N24 = 1'b0; N27 = 1'b1; N30 = 1'b0; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b0; N47 = 1'b0; N50 = 1'b1; N53 = 1'b1; N56 = 1'b1; N60 = 1'b0; N63 = 1'b1; N66 = 1'b1; N69 = 1'b1; N73 = 1'b1; N76 = 1'b1; N79 = 1'b1; N82 = 1'b0; N86 = 1'b0; N89 = 1'b0; N92 = 1'b1; N95 = 1'b0; N99 = 1'b0; N102 = 1'b1; N105 = 1'b1; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b0; N11 = 1'b0; N14 = 1'b0; N17 = 1'b1; N21 = 1'b0; N24 = 1'b1; N27 = 1'b1; N30 = 1'b0; N34 = 1'b1; N37 = 1'b0; N40 = 1'b1; N43 = 1'b1; N47 = 1'b1; N50 = 1'b1; N53 = 1'b1; N56 = 1'b1; N60 = 1'b0; N63 = 1'b1; N66 = 1'b0; N69 = 1'b0; N73 = 1'b0; N76 = 1'b0; N79 = 1'b1; N82 = 1'b0; N86 = 1'b1; N89 = 1'b0; N92 = 1'b1; N95 = 1'b0; N99 = 1'b0; N102 = 1'b1; N105 = 1'b1; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b1; N11 = 1'b0; N14 = 1'b0; N17 = 1'b1; N21 = 1'b0; N24 = 1'b0; N27 = 1'b0; N30 = 1'b1; N34 = 1'b1; N37 = 1'b0; N40 = 1'b0; N43 = 1'b1; N47 = 1'b0; N50 = 1'b0; N53 = 1'b1; N56 = 1'b1; N60 = 1'b1; N63 = 1'b0; N66 = 1'b1; N69 = 1'b1; N73 = 1'b0; N76 = 1'b1; N79 = 1'b1; N82 = 1'b0; N86 = 1'b0; N89 = 1'b1; N92 = 1'b1; N95 = 1'b1; N99 = 1'b1; N102 = 1'b1; N105 = 1'b1; N108 = 1'b0; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b1; N8 = 1'b0; N11 = 1'b0; N14 = 1'b1; N17 = 1'b1; N21 = 1'b1; N24 = 1'b0; N27 = 1'b1; N30 = 1'b0; N34 = 1'b0; N37 = 1'b1; N40 = 1'b1; N43 = 1'b1; N47 = 1'b1; N50 = 1'b0; N53 = 1'b1; N56 = 1'b1; N60 = 1'b0; N63 = 1'b1; N66 = 1'b1; N69 = 1'b1; N73 = 1'b1; N76 = 1'b1; N79 = 1'b0; N82 = 1'b1; N86 = 1'b0; N89 = 1'b0; N92 = 1'b0; N95 = 1'b0; N99 = 1'b0; N102 = 1'b1; N105 = 1'b1; N108 = 1'b1; N112 = 1'b0; N115 = 1'b0; 
#10 N1 = 1'b1; N4 = 1'b0; N8 = 1'b1; N11 = 1'b1; N14 = 1'b1; N17 = 1'b0; N21 = 1'b0; N24 = 1'b1; N27 = 1'b1; N30 = 1'b0; N34 = 1'b0; N37 = 1'b0; N40 = 1'b1; N43 = 1'b0; N47 = 1'b0; N50 = 1'b1; N53 = 1'b1; N56 = 1'b0; N60 = 1'b1; N63 = 1'b1; N66 = 1'b0; N69 = 1'b1; N73 = 1'b1; N76 = 1'b1; N79 = 1'b1; N82 = 1'b1; N86 = 1'b0; N89 = 1'b1; N92 = 1'b0; N95 = 1'b0; N99 = 1'b1; N102 = 1'b1; N105 = 1'b1; N108 = 1'b1; N112 = 1'b1; N115 = 1'b0; 
#10 N1 = 1'b0; N4 = 1'b1; N8 = 1'b0; N11 = 1'b0; N14 = 1'b0; N17 = 1'b1; N21 = 1'b0; N24 = 1'b0; N27 = 1'b1; N30 = 1'b0; N34 = 1'b1; N37 = 1'b1; N40 = 1'b0; N43 = 1'b1; N47 = 1'b0; N50 = 1'b0; N53 = 1'b1; N56 = 1'b0; N60 = 1'b1; N63 = 1'b0; N66 = 1'b1; N69 = 1'b1; N73 = 1'b1; N76 = 1'b1; N79 = 1'b1; N82 = 1'b0; N86 = 1'b1; N89 = 1'b0; N92 = 1'b1; N95 = 1'b0; N99 = 1'b1; N102 = 1'b1; N105 = 1'b0; N108 = 1'b0; N112 = 1'b1; N115 = 1'b0; 

end
endmodule
